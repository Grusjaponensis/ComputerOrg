module StallController();
    
endmodule //StallController
