module led(
    input [3:0] x,
    output a, b, c, d, e, f, g
);
    assign a = (~x[0] & x[3]) | (~x[0] & x[2]) | (x[0] & ~x[1] & ~x[2]) | (x[0] & ~x[3]) | (x[1] & x[2]);
    assign b = (~x[2] & ~x[3]) | (x[2] & ~x[3]) | (x[0] & x[2]) | (x[0] & x[1]);
    assign c = (~x[1] & ~x[3]) | (x[2] & ~x[3]) | (x[0] & x[2]) | (x[0] & x[1]);
    assign d = (x[1] & ~x[2] & x[3]) | (~x[0] & ~x[1] & ~x[3]) | (~x[0] & ~x[1] & x[2]) | (~x[0] & x[2] & ~x[3]) | (~x[1] & ~x[2] & ~x[3]) | (x[0] & ~x[2]) | (~x[1] & x[2] & x[3]) | (x[1] & x[2] & ~x[3]);
    assign e = ~x[0] | ~x[1] | (x[2] & x[3]);
    assign f = (x[0] & ~x[2] & ~x[3]) | (~x[0] & x[2] & x[3]) | (x[0] & ~x[1] & ~x[3]) | (x[0] & ~x[2] & x[3]) | (~x[0] & ~x[1] & x[3]);
    assign g = (~x[1] & x[2]) | (x[0] & ~x[1]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & x[1] & ~x[3]) | (x[1] & ~x[2] & x[3]) | (x[2] & ~x[3]) | (x[0] & x[3]);
endmodule