module ForwardController();
    
endmodule //ForwardController
