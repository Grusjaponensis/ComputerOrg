`timescale 1ns / 1ps
module intcheck_tb;

	// Inputs
	reg clk;
	reg reset;
	reg [7:0] in;

	// Outputs
	wire out;

	// Instantiate the Unit Under Test (UUT)
	intcheck uut (
		.clk(clk), 
		.reset(reset), 
		.in(in), 
		.out(out)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		in = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		// #2;
        // in = " ";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "a";
        // #2;
        // in = ";";
        // #2;
        // in = " ";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = ";";

        // #2;
        // in = " ";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "a";
        // #2;
        // in = "_";
        // #2;
        // in = ",";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "p";
        // #2;
        // in = ";";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = ";";

        // #2;
        // in = " ";
        // #2;
        // in = " ";
        // #2;
        // in = "\t";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "\t";
        // #2;
        // in = "9";
        // #2;
        // in = "n";
        // #2;
        // in = "p";
        // #2;
        // in = " ";
        // #2;
        // in = ";";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = "a";
        // #2;
        // in = "_";
        // #2;
        // in = ",";
        // #2;
        // in = ";";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "p";
        // #2;
        // in = ";";

        // #2;
        // in = " ";
        // #2;
        // in = " ";
        // #2;
        // in = "\t";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        // in = ";";
        // #2;
        // in = ";";
        // #2;
        // in = "i";
        // #2;
        // in = "n";
        // #2;
        // in = "t";
        // #2;
        // in = " ";
        // #2;
        in = "i";
        #2;
        in = "n";
        #2;
        in = "t";
        #2;
        in = " ";
        #2;
        in = "a";
        #2;
        in = " ";
        #2;
        in = "B";
        #2;
        in = ";";
        #2;
        in = "1";
        #2;
        in = ",";
        #2;
        in = " ";
        #2;
        in = "i";
        #2;
        in = "n";
        #2;
        in = "p";
        #2;
        in = "_";
        #2;
        in = "3";
        #2;
        in = " ";
        #2;
        in = ",";
        #2;
        in = " ";
        #2;
        in = "\t";
        #2;
        in = "9";
        #2;
        in = "0";
        #2;
        in = "a";
        #2;
        in = ";";
        #2;
        in = "i";
        #2;
        in = "n";
        #2;
        in = "t";
        #2;
        in = " ";
        #2;
        #2;
        in = "d";
        #2;
        in = ",";
        #2;
        in = "_";
        #2;
        in = "9";
        #2;
        in = ";";
        #2;
        in = "i";
        #2;
        in = "n";
        #2;
        in = "t";
        #2;
        in = " ";
        #2;
        in = "i";
        #2;
        in = "n";
        #2;
        in = "t";
        #2;
        in = ";";
	end
    always #1 clk = ~clk;
endmodule